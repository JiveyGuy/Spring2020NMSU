library IEEE;
use 	IEEE.STD_Logic_1164.All;
use 	IEEE.NUMERIC_STD.All;

Library EE_212_ALU;
use 	EE_212_ALU.ALU.all;

Library EE_212_NIAG;
use 	EE_212_NIAG.NIAG.all;

ENTITY NIAG IS 

	PORT( 
		Target	:	IN	STD_LOGIC_VECTOR(25 DOWNTO 0);
		Immed	:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		Reg	:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		Xshft	:	IN	STD_LOGIC;
		PCin	:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		Cond	:	IN	STD_LOGIC_VECTOR(2 DOWNTO 0);
		Sel	:	IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		Stat	:	IN	STAT_SIGNL_REC;
		MemAdrs	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
		RtnAdrs	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEHAVIORAL OF NIAG IS 
		
SIGNAL NSA 	 : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL AbsltAdrs : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL RegAdrs   : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL RelAdrs   : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL RetAdrs   : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN 
	FOO : NIAG_NSA   PORT MAP( PCin, NSA);
	FO1 : NIAG_Abslt PORT MAP( Target, NSA, AbsltAdrs);
	FO2 : NIAG_Reg   PORT MAP( Reg, Regadrs );
	FO3 : NIAG_Rel   PORT MAP( Immed, XShft, NSA, RelAdrs );
	FO4 : NIAG_Rtn   PORT MAP( PCin, RtnAdrs );
	FO5 : NIAG_Mux   PORT MAP( NSA, AbsltAdrs, RelAdrs, RegAdrs, Cond, Sel, Stat, MemAdrs);
END ARCHITECTURE;