library IEEE;
use 	IEEE.STD_Logic_1164.All;
use 	IEEE.NUMERIC_STD.All;

Library EE_212_ALU;
use 	EE_212_ALU.ALU.all;

Library EE_212_DECODER;
use 	EE_212_DECODER.DecodeLogic.all;

ENTITY NIAG_Rtn IS 
	PORT(	PC	:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		RtnAdrs	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF NIAG_Rtn IS 
	BEGIN PROCESS ( PC ) BEGIN
		RtnAdrs <= STD_LOGIC_VECTOR(Unsigned(PC) + 8);
	END PROCESS;
END ARCHITECTURE;

-- This just gives Reg to RegAdrs
